

 
 
 




window new WaveWindow  -name  "Waves for BMG Example Design"
waveform  using  "Waves for BMG Example Design"

      waveform add -signals /downtube_tb/status
      waveform add -signals /downtube_tb/downtube_synth_inst/bmg_port/CLKA
      waveform add -signals /downtube_tb/downtube_synth_inst/bmg_port/ADDRA
      waveform add -signals /downtube_tb/downtube_synth_inst/bmg_port/DOUTA

console submit -using simulator -wait no "run"
