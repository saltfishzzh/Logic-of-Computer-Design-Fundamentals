`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    17:40:53 12/10/2014 
// Design Name: 
// Module Name:    prom_DMH 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module prom_DMH(
input wire [3:0] addr,
output wire [0:31] M
    );
	 reg[0:31] rom[0:15];
	 parameter data = {
				32'b000000001111111111111111000000,
				32'b000000000000000000000000000000,
				32'b000000000000000000000001110000,
				32'b100000000000000000000000000000,
				32'b100000000000000000000000000000,
				32'b100000000000000000000000000000,
				32'b000000001110000000011100000000,
				32'b000000000000000000000000000000,
				32'b000000000000000000000000000000,
				32'b000000000000000000000000000000,
				32'b000000000000111000000000000000,
				32'b000000000000000000000000000001,
				32'b000000000000000000000000000001,
				32'b000000111000000000000000000001,
				32'b000000000000000000000000000000,
				32'b000000000000000000001100000000 };
		integer i;
		initial 
		begin
			for(i = 0; i < 16; i = i + 1)
				rom[i] = data[(511-32*i)-:32];
		end

		assign M = rom[addr];

endmodule
