`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    20:17:55 01/11/2015 
// Design Name: 
// Module Name:    CountScore 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module CountScore(
input wire clk,
input wire[7:0] score,
input wire[5:0] rom1_addr,
input wire[5:0] rom2_addr,
output wire[0:31] M1,
output wire[0:31] M2
    );
	 
parameter data0={
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111100000000001111111111,
32'b11111111110000000000000011111111,
32'b11111111100000000000000000111111,
32'b11111111000000000000000000011111,
32'b11111110000000011110000000001111,
32'b11111100000000111111000000001111,
32'b11111100000001111111100000000111,
32'b11111000000011111111110000000111,
32'b11110000000011111111110000000011,
32'b11110000000011111111110000000011,
32'b11100000000111111111111000000011,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000001,
32'b11100000000111111111111000000011,
32'b11100000000111111111111000000011,
32'b11110000000111111111111000000011,
32'b11110000000011111111111000000011,
32'b11111000000001111111110000000111,
32'b11111100000000111111100000001111,
32'b11111110000000011110000000001111,
32'b11111111000000000000000000011111,
32'b11111111100000000000000000111111,
32'b11111111110000000000000011111111,
32'b11111111111100000000001111111111,
32'b11111111111111111111111111111111
};
parameter data1={
32'b11111111111111111111111111111111,
32'b11111111111111100000000000001111,
32'b11111111111110000000000000001111,
32'b11111111111000000000000000001111,
32'b11111111000000000000000000001111,
32'b11111000000000000000000000001111,
32'b10000000000000000000000000001111,
32'b10000000000000000000000000001111,
32'b10000000000000000000000000001111,
32'b10000000000011100000000000000111,
32'b10000000011111100000000000001111,
32'b10000011111111100000000000001111,
32'b10111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111100000000000001111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};
parameter data2={
32'b11111111111111111111111111111111,
32'b11111111111000000000011111111111,
32'b11111111000000000000000011111111,
32'b11111100000000000000000000111111,
32'b11111000000000000000000000011111,
32'b11110000000000011000000000001111,
32'b11110000000001111111000000001111,
32'b11100000000011111111100000000111,
32'b11100000000111111111100000000111,
32'b11100000000111111111100000000111,
32'b11100000000111111111110000000011,
32'b11111111111111111111110000000011,
32'b11111111111111111111100000000111,
32'b11111111111111111111100000000111,
32'b11111111111111111111000000000111,
32'b11111111111111111111000000001111,
32'b11111111111111111110000000001111,
32'b11111111111111111100000000011111,
32'b11111111111111111000000000111111,
32'b11111111111111110000000001111111,
32'b11111111111111100000000001111111,
32'b11111111111111000000000011111111,
32'b11111111111110000000001111111111,
32'b11111111111100000000001111111111,
32'b11111111111000000000111111111111,
32'b11111111100000000001111111111111,
32'b11111111000000000011111111111111,
32'b11111110000000000111111111111111,
32'b11111100000000001111111111111111,
32'b11110000000000111111111111111111,
32'b11100000000001111111111111111111,
32'b11000000000011111111111111111111,
32'b11000000001111111111111111111111,
32'b11000000001111111111111111111111,
32'b11000000000000000000000000000011,
32'b11000000000000000000000000000011,
32'b11000000000000000000000000000011,
32'b11000000000000000000000000000011,
32'b11000000000000000000000000000011,
32'b11111111111111111111111111111111
};
parameter data3={
32'b11111111111111111111111111111111,
32'b11111111111000000000011111111111,
32'b11111111100000000000000011111111,
32'b11111110000000000000000000111111,
32'b11111100000000000000000000011111,
32'b11111100000000001110000000001111,
32'b11111000000000111111000000001111,
32'b11111000000001111111100000000111,
32'b11110000000011111111110000000111,
32'b11110000000011111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111100000000111,
32'b11111111111111111111100000001111,
32'b11111111111111111111000000011111,
32'b11111111111111111100000000111111,
32'b11111111111100000000000001111111,
32'b11111111111110000000001111111111,
32'b11111111111110000000001111111111,
32'b11111111111110000000000011111111,
32'b11111111111110000000000000111111,
32'b11111111111111111100000000111111,
32'b11111111111111111111000000001111,
32'b11111111111111111111100000001111,
32'b11111111111111111111100000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11110000000111111111110000000111,
32'b11110000000111111111110000000111,
32'b11110000000011111111100000000111,
32'b11110000000011111111100000000111,
32'b11111000000000111111000000001111,
32'b11111000000000001100000000011111,
32'b11111100000000000000000000111111,
32'b11111110000000000000000001111111,
32'b11111111100000000000001111111111,
32'b11111111111111000111111111111111,
32'b11111111111111111111111111111111
};
parameter data4={
32'b11111111111111111111111111111111,
32'b11111111111111111000000011111111,
32'b11111111111111110000000011111111,
32'b11111111111111110000000011111111,
32'b11111111111111100000000011111111,
32'b11111111111111000000000011111111,
32'b11111111111111000000000011111111,
32'b11111111111110000000000011111111,
32'b11111111111100000000000011111111,
32'b11111111111000000000000011111111,
32'b11111111111000000100000011111111,
32'b11111111110000001100000011111111,
32'b11111111110000011100000011111111,
32'b11111111100000111100000011111111,
32'b11111111000000111100000011111111,
32'b11111110000001111100000011111111,
32'b11111110000011111100000011111111,
32'b11111100000111111100000011111111,
32'b11111000000111111100000011111111,
32'b11111000001111111100000011111111,
32'b11110000011111111100000011111111,
32'b11100000111111111100000011111111,
32'b11000001111111111100000011111111,
32'b11000001111111111100000011111111,
32'b11000001111111111100000011111111,
32'b11000000000000000000000000000011,
32'b11000000000000000000000000000011,
32'b11000000000000000000000000000011,
32'b11000000000000000000000000000011,
32'b11000000000000000000000000000011,
32'b11111111111111111100000011111111,
32'b11111111111111111100000011111111,
32'b11111111111111111100000001111111,
32'b11111111111111111100000001111111,
32'b11111111111111111100000001111111,
32'b11111111111111111100000001111111,
32'b11111111111111111100000001111111,
32'b11111111111111111100000001111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};
parameter data5={
32'b11111111111111111111111111111111,
32'b11110000000000000000000000011111,
32'b11110000000000000000000000011111,
32'b11110000000000000000000000011111,
32'b11110000000000000000000000011111,
32'b11110000001111111111111111111111,
32'b11110000001111111111111111111111,
32'b11110000001111111111111111111111,
32'b11110000001111111111111111111111,
32'b11110000001111111111111111111111,
32'b11110000001111111111111111111111,
32'b11110000001111111111111111111111,
32'b11110000001111111111111111111111,
32'b11110000001111111111111111111111,
32'b11110000001111000000001111111111,
32'b11110000001100000000000001111111,
32'b11110000000000000000000000111111,
32'b11110000000000000000000000011111,
32'b11110000000000011100000000011111,
32'b11110000000001111110000000001111,
32'b11110000000011111111000000001111,
32'b11110000000111111111100000001111,
32'b11111111111111111111110000001111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11110000000111111111100000001111,
32'b11110000000111111111100000001111,
32'b11110000000011111111000000011111,
32'b11111000000001111100000000011111,
32'b11111000000000000000000000111111,
32'b11111100000000000000000001111111,
32'b11111111000000000000000111111111,
32'b11111111110000000000111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111
};
parameter data6={
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111111111110001111111111111,
32'b11111111111000000000000011111111,
32'b11111111100000000000000000111111,
32'b11111110000000000000000000001111,
32'b11111100000000000000000000000111,
32'b11111100000000111111000000000111,
32'b11111000000001111111100000000011,
32'b11110000000011111111110000000011,
32'b11110000000111111111110000000011,
32'b11100000000111111111111111111111,
32'b11100000000111111111111111111111,
32'b11100000001111111111111111111111,
32'b11100000001111111111111111111111,
32'b11000000001111111111111111111111,
32'b11000000001111110000011111111111,
32'b11000000001110000000000001111111,
32'b11000000001000000000000000011111,
32'b11000000000000000000000000001111,
32'b11000000000000001000000000000111,
32'b11000000000001111111000000000011,
32'b11000000000011111111100000000011,
32'b11000000000011111111110000000011,
32'b11000000000111111111110000000001,
32'b11000000001111111111111000000001,
32'b11000000001111111111111000000001,
32'b11000000001111111111111000000001,
32'b11000000001111111111111000000001,
32'b11000000001111111111111000000001,
32'b11000000001111111111110000000001,
32'b11000000000111111111110000000001,
32'b11000000000111111111110000000011,
32'b11100000000011111111100000000011,
32'b11110000000001111111000000000111,
32'b11111000000000001000000000001111,
32'b11111100000000000000000000011111,
32'b11111110000000000000000011111111,
32'b11111111000000000000000111111111,
32'b11111111111111111111111111111111
};
parameter data7={
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11100000000000000000000000000011,
32'b11100000000000000000000000000011,
32'b11100000000000000000000000000011,
32'b11100000000000000000000000000011,
32'b11100000000000000000000000000011,
32'b11111111111111111111111000000011,
32'b11111111111111111111110000000011,
32'b11111111111111111111110000000011,
32'b11111111111111111111100000000111,
32'b11111111111111111111100000000111,
32'b11111111111111111111000000000111,
32'b11111111111111111111000000001111,
32'b11111111111111111111000000001111,
32'b11111111111111111110000000011111,
32'b11111111111111111110000000011111,
32'b11111111111111111100000000111111,
32'b11111111111111111100000000111111,
32'b11111111111111111000000001111111,
32'b11111111111111111000000001111111,
32'b11111111111111110000000001111111,
32'b11111111111111110000000011111111,
32'b11111111111111100000000011111111,
32'b11111111111111100000000111111111,
32'b11111111111111000000000111111111,
32'b11111111111111000000001111111111,
32'b11111111111111000000001111111111,
32'b11111111111110000000011111111111,
32'b11111111111110000000011111111111,
32'b11111111111100000000111111111111,
32'b11111111111100000000111111111111,
32'b11111111111000000000111111111111,
32'b11111111111000000001111111111111,
32'b11111111110000000001111111111111,
32'b11111111110000000011111111111111,
32'b11111111110000000111111111111111,
32'b11111111100000000111111111111111,
32'b11111111000000001111111111111111,
32'b11111111111111111111111111111111
};
parameter data8={
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111110000000000001111111111,
32'b11111111000000000000000011111111,
32'b11111110000000000000000000111111,
32'b11111100000000000000000000011111,
32'b11111000000001111100000000011111,
32'b11110000000011111111000000001111,
32'b11110000000111111111100000001111,
32'b11110000001111111111110000001111,
32'b11110000001111111111110000000111,
32'b11110000001111111111110000000111,
32'b11110000001111111111110000001111,
32'b11110000001111111111110000001111,
32'b11110000000111111111100000001111,
32'b11111000000011111111000000011111,
32'b11111000000001111110000000111111,
32'b11111110001000000000000001111111,
32'b11111111100000000000001111111111,
32'b11111111110000000000001111111111,
32'b11111111110000000000001111111111,
32'b11111110000000000000001001111111,
32'b11111100000000011000000000111111,
32'b11111000000011111111000000011111,
32'b11110000000111111111000000011111,
32'b11110000000111111111100000000111,
32'b11100000001111111111110000000111,
32'b11100000001111111111110000000111,
32'b11100000001111111111110000000111,
32'b11100000001111111111110000000111,
32'b11100000001111111111110000000111,
32'b11100000001111111111110000000111,
32'b11100000000111111111100000001111,
32'b11110000000111111111000000001111,
32'b11110000000011111110000000011111,
32'b11111000000000011000000000011111,
32'b11111100000000000000000000111111,
32'b11111110000000000000000011111111,
32'b11111111110000000000001111111111,
32'b11111111111111111111111111111111
};
parameter data9={
32'b11111111111111111111111111111111,
32'b11111111111111111111111111111111,
32'b11111111110000000000001111111111,
32'b11111111000000000000000011111111,
32'b11111110000000000000000000111111,
32'b11111000000000000000000000011111,
32'b11110000000000111110000000001111,
32'b11110000000011111111000000001111,
32'b11100000000111111111100000000111,
32'b11100000000111111111110000000111,
32'b11100000001111111111110000000011,
32'b11000000001111111111111000000011,
32'b11000000001111111111111000000011,
32'b11000000001111111111111000000011,
32'b11000000001111111111111000000011,
32'b11000000001111111111110000000011,
32'b11100000001111111111110000000011,
32'b11100000000111111111110000000011,
32'b11100000000011111111100000000011,
32'b11110000000000111110000000000011,
32'b11111000000000000000000000000011,
32'b11111100000000000000000000000011,
32'b11111110000000000000000000000011,
32'b11111111100000000000111000000011,
32'b11111111111110001111111000000011,
32'b11111111111111111111111000000011,
32'b11111111111111111111111000000011,
32'b11111111111111111111111000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11111111111111111111110000000111,
32'b11100000000111111111100000000111,
32'b11100000000111111111100000001111,
32'b11100000000011111111000000001111,
32'b11110000000001111110000000011111,
32'b11110000000000000000000000111111,
32'b11111000000000000000000001111111,
32'b11111110000000000000000011111111,
32'b11111111100000000000011111111111,
32'b11111111111111111111111111111111
};

reg[0:31] rom1[0:39];
reg[0:31] rom2[0:39];
integer i;

always@(posedge clk) begin
	case(score[7:4])
	0:for(i=0;i<40;i=i+1) rom1[i] = data0[(1279-32*i)-:32];
	1:for(i=0;i<40;i=i+1) rom1[i] = data1[(1279-32*i)-:32];
	2:for(i=0;i<40;i=i+1) rom1[i] = data2[(1279-32*i)-:32];
	3:for(i=0;i<40;i=i+1) rom1[i] = data3[(1279-32*i)-:32];
	4:for(i=0;i<40;i=i+1) rom1[i] = data4[(1279-32*i)-:32];
	5:for(i=0;i<40;i=i+1) rom1[i] = data5[(1279-32*i)-:32];
	6:for(i=0;i<40;i=i+1) rom1[i] = data6[(1279-32*i)-:32];
	7:for(i=0;i<40;i=i+1) rom1[i] = data7[(1279-32*i)-:32];
	8:for(i=0;i<40;i=i+1) rom1[i] = data8[(1279-32*i)-:32];
	default:for(i=0;i<40;i=i+1) rom1[i] = data9[(1279-32*i)-:32];
	endcase//endcase for score[7:4]
	case(score[3:0])
	0:for(i=0;i<40;i=i+1) rom2[i] = data0[(1279-32*i)-:32];
	1:for(i=0;i<40;i=i+1) rom2[i] = data1[(1279-32*i)-:32];
	2:for(i=0;i<40;i=i+1) rom2[i] = data2[(1279-32*i)-:32];
	3:for(i=0;i<40;i=i+1) rom2[i] = data3[(1279-32*i)-:32];
	4:for(i=0;i<40;i=i+1) rom2[i] = data4[(1279-32*i)-:32];
	5:for(i=0;i<40;i=i+1) rom2[i] = data5[(1279-32*i)-:32];
	6:for(i=0;i<40;i=i+1) rom2[i] = data6[(1279-32*i)-:32];
	7:for(i=0;i<40;i=i+1) rom2[i] = data7[(1279-32*i)-:32];
	8:for(i=0;i<40;i=i+1) rom2[i] = data8[(1279-32*i)-:32];
	default:for(i=0;i<40;i=i+1) rom2[i] = data9[(1279-32*i)-:32];
	endcase//endcase for score[3:0]
end

assign M1 = rom1[rom1_addr];
assign M2 = rom2[rom2_addr];

endmodule
